`timescale 1ns / 10ps

module % #(
    // parameters
) (
    input clk, n_rst
);



endmodule

