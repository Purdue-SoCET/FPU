module decoder (

);

endmodule
